component highlevel.ServerKettle

endpoints {
    service : highlevel.ServiceKettle
}
