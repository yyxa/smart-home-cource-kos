component highlevel.ServerChecker

endpoints {
    service : highlevel.ServiceChecker
}
