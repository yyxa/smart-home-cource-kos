component highlevel.ServerKeys

endpoints {
    service : highlevel.ServiceKeys
}
